// char gaussian_bit_pattern_31_x_a[256] = { 8,4,-11,7,2,1,-2,-13,-13,10,-13,-11,7,-4,-13,-9,12,-3,-6,11,4,5,3,-8,-2,-13,-7,-4,-10,5,5,1,9,4,2,-4,-8,4,0,-13,-3,-6,8,0,7,-13,10,-6,10,-13,-13,3,5,-1,3,2,-13,-13,-13,-7,6,-9,-2,-12,3,-7,-3,2,-11,-1,5,-4,-9,-12,10,7,-7,-4,7,-7,-13,-3,7,-13,1,2,-4,-1,7,1,9,-1,-13,7,12,6,5,2,3,2,9,-8,-11,1,6,2,6,3,7,-11,-10,-5,-10,8,4,-10,4,-2,-5,7,-9,-5,8,-9,1,7,-2,11,-12,3,5,0,-9,0,-1,5,3,-13,-5,-4,6,-7,-13,1,4,-2,2,-2,4,-6,-3,7,4,-13,7,7,-7,-8,-13,2,10,-6,8,2,-11,-12,-11,5,-2,-1,-13,-10,-3,2,-9,-4,-4,-6,6,-13,11,7,-1,-4,-7,-13,-7,-8,-5,-13,1,1,9,5,-1,-9,-1,-13,8,2,7,-10,-10,4,3,-4,5,4,-9,0,-12,3,-10,8,-8,2,10,6,-7,-3,-1,-3,-8,4,2,6,3,11,-3,4,2,-10,-13,-13,6,0,-13,-9,-13,5,2,-1,9,11,3,-1,3,-13,5,8,7,-10,7,9,7,-1};
// char gaussian_bit_pattern_31_y_a[256] = {-3,2,9,-12,-13,-7,-10,-13,-3,4,-8,7,7,-5,2,0,-6,6,-13,-13,7,-3,-7,-7,11,12,3,2,-12,-12,-6,0,11,7,-1,-12,-5,11,-8,-2,-2,9,12,9,-5,-6,7,-3,-9,8,0,3,7,7,-10,-4,0,-7,3,12,-10,-1,-5,5,-10,-7,-2,9,-13,6,-3,-13,-6,-10,2,12,-13,9,-1,6,11,7,-8,-7,-3,-6,3,-13,1,-1,1,-9,-13,7,-5,3,-13,-12,8,6,-12,4,12,12,-9,3,3,-3,8,-5,11,-8,5,-1,-6,12,-2,0,-8,-6,-13,-13,-8,-11,-8,-4,1,-6,-9,7,5,-4,12,7,2,11,5,-4,9,-7,5,6,6,-10,1,-2,-12,-13,1,-10,-13,5,-2,9,1,-8,-4,11,6,4,-5,-5,-3,-12,-2,-13,0,-3,-13,-8,-11,-2,9,-3,-13,6,12,-11,-3,11,11,-5,12,-8,1,-12,-2,5,-1,7,5,0,12,-8,11,-3,-10,1,-11,-13,-13,-10,-8,-6,12,2,-13,-13,9,3,1,2,-10,-13,-12,2,6,8,10,-9,-13,-7,-2,2,-5,-9,-1,-1,0,-11,-4,-6,7,12,0,-1,3,8,-6,-9,7,-6,5,-3,0,4,-6,0,8,9,-4,4,3,-7,0,-6};
// char gaussian_bit_pattern_31_x_b[256] = {9,7,-8,12,2,1,-2,-11,-12,11,-8,-9,12,-3,-12,-7,12,-2,-4,12,5,10,6,-6,-1,-8,-5,-3,-6,6,7,4,11,4,4,-2,-7,9,1,-8,-2,-4,10,1,11,-11,12,-6,12,-8,-8,7,10,1,5,3,-13,-12,-11,-4,12,-7,0,-7,8,-4,-1,5,-5,0,5,-4,-9,-8,12,12,-6,-3,12,-5,-12,-2,12,-11,12,3,-2,1,8,3,12,-1,-10,10,12,7,6,2,4,12,10,-7,-4,2,7,3,11,8,9,-6,-5,-3,-9,12,6,-8,6,-2,-5,10,-8,-5,9,-9,1,9,-1,12,-6,7,10,2,-5,2,1,7,6,-8,-3,-3,8,-6,-5,3,8,2,12,0,9,-3,-1,12,5,-9,8,7,-7,-7,-12,3,12,-6,9,2,-10,-7,-10,11,-1,0,-12,-10,-2,3,-4,-3,-2,-4,6,-5,12,12,0,-3,-6,-8,-6,-6,-4,-8,5,10,10,10,1,-6,1,-8,10,3,12,-5,-8,8,8,-3,10,5,-4,3,-6,4,-10,12,-6,3,11,8,-6,-3,-1,-3,-8,12,3,11,7,12,-3,4,2,-8,-11,-11,11,1,-9,-6,-8,8,3,-1,11,12,3,0,4,-10,12,9,8,-10,12,10,12,0};
// char gaussian_bit_pattern_31_y_b[256] = {5,-12,2,-13,12,6,-4,-8,-9,9,-9,12,6,0,-3,5,-1,12,-8,-8,1,-3,12,-2,-10,10,-3,7,11,-7,-1,-5,-13,12,4,7,-10,12,-13,2,3,-9,7,3,-10,0,1,12,-4,-12,-4,8,-7,-12,6,-10,5,12,8,7,8,-6,12,5,-13,5,-7,-11,-13,-1,2,12,6,-4,-3,12,5,4,2,1,5,-6,-7,-12,12,0,-13,9,-6,12,6,3,5,12,9,11,10,3,-6,-13,3,9,-6,-8,-4,-2,0,-8,3,-4,10,12,0,-6,-11,7,7,12,2,12,-8,-2,-13,0,-2,1,-4,-11,4,12,8,8,-13,12,7,-9,-8,9,-3,-12,0,12,-2,10,-4,-13,12,-6,3,-5,1,-11,-7,-5,6,6,1,-8,-8,9,3,7,-8,8,3,-9,-5,8,12,9,-5,11,-13,2,0,-10,-7,9,11,5,6,-2,7,-2,7,-13,-8,-9,5,10,-13,-13,-1,-9,-13,2,12,-10,-6,-6,-9,-7,-13,5,-13,-3,-12,-1,3,-9,1,-8,9,12,-5,7,-8,-12,5,9,5,4,3,12,11,-13,12,4,6,12,1,1,1,-13,-13,4,-2,-3,-2,10,-9,-1,-2,-8,5,10,5,5,11,-6,-12,9,4,-2,-2,-11};

// float cos_angle = std::cos(orientation);
// float sin_angle = std::sin(orientation);

// x1 = round((gaussian_bit_pattern_31_x_a[index]*cos_angle - gaussian_bit_pattern_31_y_a[index]*sin_angle));
// y1 = round((gaussian_bit_pattern_31_x_a[index]*sin_angle + gaussian_bit_pattern_31_y_a[index]*cos_angle));
// x2 = round((gaussian_bit_pattern_31_x_b[index]*cos_angle - gaussian_bit_pattern_31_y_b[index]*sin_angle));
// y2 = round((gaussian_bit_pattern_31_x_b[index]*sin_angle + gaussian_bit_pattern_31_y_b[index]*cos_angle));

module LUT
(
    input [7:0] i_num,
    output logic [7:0] o_xa,
    output logic [7:0] o_ya,
    output logic [7:0] o_xb,
    output logic [7:0] o_yb
);

    always_comb begin
        case(i_num)
            0: begin
                o_xa = 8'd8;
                o_ya = -8'd3;
                o_xb = 8'd9;
                o_yb = 8'd5;
            end
            1: begin
                o_xa = 8'd4;
                o_ya = 8'd2;
                o_xb = 8'd7;
                o_yb = -8'd12;
            end
            2: begin
                o_xa = -8'd11;
                o_ya = 8'd9;
                o_xb = -8'd8;
                o_yb = 8'd2;
            end
            3: begin
                o_xa = 8'd7;
                o_ya = -8'd12;
                o_xb = 8'd12;
                o_yb = -8'd13;
            end
            4: begin
                o_xa = 8'd2;
                o_ya = -8'd13;
                o_xb = 8'd2;
                o_yb = 8'd12;
            end
            5: begin
                o_xa = 8'd1;
                o_ya = -8'd7;
                o_xb = 8'd1;
                o_yb = 8'd6;
            end
            6: begin
                o_xa = -8'd2;
                o_ya = -8'd10;
                o_xb = -8'd2;
                o_yb = -8'd4;
            end
            7: begin
                o_xa = -8'd13;
                o_ya = -8'd13;
                o_xb = -8'd11;
                o_yb = -8'd8;
            end
            8: begin
                o_xa = -8'd13;
                o_ya = -8'd3;
                o_xb = -8'd12;
                o_yb = -8'd9;
            end
            9: begin
                o_xa = 8'd10;
                o_ya = 8'd4;
                o_xb = 8'd11;
                o_yb = 8'd9;
            end
            10: begin
                o_xa = -8'd13;
                o_ya = -8'd8;
                o_xb = -8'd8;
                o_yb = -8'd9;
            end
            11: begin
                o_xa = -8'd11;
                o_ya = 8'd7;
                o_xb = -8'd9;
                o_yb = 8'd12;
            end
            12: begin
                o_xa = 8'd7;
                o_ya = 8'd7;
                o_xb = 8'd12;
                o_yb = 8'd6;
            end
            13: begin
                o_xa = -8'd4;
                o_ya = -8'd5;
                o_xb = -8'd3;
                o_yb = 8'd0;
            end
            14: begin
                o_xa = -8'd13;
                o_ya = 8'd2;
                o_xb = -8'd12;
                o_yb = -8'd3;
            end
            15: begin
                o_xa = -8'd9;
                o_ya = 8'd0;
                o_xb = -8'd7;
                o_yb = 8'd5;
            end
            16: begin
                o_xa = 8'd12;
                o_ya = -8'd6;
                o_xb = 8'd12;
                o_yb = -8'd1;
            end
            17: begin
                o_xa = -8'd3;
                o_ya = 8'd6;
                o_xb = -8'd2;
                o_yb = 8'd12;
            end
            18: begin
                o_xa = -8'd6;
                o_ya = -8'd13;
                o_xb = -8'd4;
                o_yb = -8'd8;
            end
            19: begin
                o_xa = 8'd11;
                o_ya = -8'd13;
                o_xb = 8'd12;
                o_yb = -8'd8;
            end
            20: begin
                o_xa = 8'd4;
                o_ya = 8'd7;
                o_xb = 8'd5;
                o_yb = 8'd1;
            end
            21: begin
                o_xa = 8'd5;
                o_ya = -8'd3;
                o_xb = 8'd10;
                o_yb = -8'd3;
            end
            22: begin
                o_xa = 8'd3;
                o_ya = -8'd7;
                o_xb = 8'd6;
                o_yb = 8'd12;
            end
            23: begin
                o_xa = -8'd8;
                o_ya = -8'd7;
                o_xb = -8'd6;
                o_yb = -8'd2;
            end
            24: begin
                o_xa = -8'd2;
                o_ya = 8'd11;
                o_xb = -8'd1;
                o_yb = -8'd10;
            end
            25: begin
                o_xa = -8'd13;
                o_ya = 8'd12;
                o_xb = -8'd8;
                o_yb = 8'd10;
            end
            26: begin
                o_xa = -8'd7;
                o_ya = 8'd3;
                o_xb = -8'd5;
                o_yb = -8'd3;
            end
            27: begin
                o_xa = -8'd4;
                o_ya = 8'd2;
                o_xb = -8'd3;
                o_yb = 8'd7;
            end
            28: begin
                o_xa = -8'd10;
                o_ya = -8'd12;
                o_xb = -8'd6;
                o_yb = 8'd11;
            end
            29: begin
                o_xa = 8'd5;
                o_ya = -8'd12;
                o_xb = 8'd6;
                o_yb = -8'd7;
            end
            30: begin
                o_xa = 8'd5;
                o_ya = -8'd6;
                o_xb = 8'd7;
                o_yb = -8'd1;
            end
            31: begin
                o_xa = 8'd1;
                o_ya = 8'd0;
                o_xb = 8'd4;
                o_yb = -8'd5;
            end
            32: begin
                o_xa = 8'd9;
                o_ya = 8'd11;
                o_xb = 8'd11;
                o_yb = -8'd13;
            end
            33: begin
                o_xa = 8'd4;
                o_ya = 8'd7;
                o_xb = 8'd4;
                o_yb = 8'd12;
            end
            34: begin
                o_xa = 8'd2;
                o_ya = -8'd1;
                o_xb = 8'd4;
                o_yb = 8'd4;
            end
            35: begin
                o_xa = -8'd4;
                o_ya = -8'd12;
                o_xb = -8'd2;
                o_yb = 8'd7;
            end
            36: begin
                o_xa = -8'd8;
                o_ya = -8'd5;
                o_xb = -8'd7;
                o_yb = -8'd10;
            end
            37: begin
                o_xa = 8'd4;
                o_ya = 8'd11;
                o_xb = 8'd9;
                o_yb = 8'd12;
            end
            38: begin
                o_xa = 8'd0;
                o_ya = -8'd8;
                o_xb = 8'd1;
                o_yb = -8'd13;
            end
            39: begin
                o_xa = -8'd13;
                o_ya = -8'd2;
                o_xb = -8'd8;
                o_yb = 8'd2;
            end
            40: begin
                o_xa = -8'd3;
                o_ya = -8'd2;
                o_xb = -8'd2;
                o_yb = 8'd3;
            end
            41: begin
                o_xa = -8'd6;
                o_ya = 8'd9;
                o_xb = -8'd4;
                o_yb = -8'd9;
            end
            42: begin
                o_xa = 8'd8;
                o_ya = 8'd12;
                o_xb = 8'd10;
                o_yb = 8'd7;
            end
            43: begin
                o_xa = 8'd0;
                o_ya = 8'd9;
                o_xb = 8'd1;
                o_yb = 8'd3;
            end
            44: begin
                o_xa = 8'd7;
                o_ya = -8'd5;
                o_xb = 8'd11;
                o_yb = -8'd10;
            end
            45: begin
                o_xa = -8'd13;
                o_ya = -8'd6;
                o_xb = -8'd11;
                o_yb = 8'd0;
            end
            46: begin
                o_xa = 8'd10;
                o_ya = 8'd7;
                o_xb = 8'd12;
                o_yb = 8'd1;
            end
            47: begin
                o_xa = -8'd6;
                o_ya = -8'd3;
                o_xb = -8'd6;
                o_yb = 8'd12;
            end
            48: begin
                o_xa = 8'd10;
                o_ya = -8'd9;
                o_xb = 8'd12;
                o_yb = -8'd4;
            end
            49: begin
                o_xa = -8'd13;
                o_ya = 8'd8;
                o_xb = -8'd8;
                o_yb = -8'd12;
            end
            50: begin
                o_xa = -8'd13;
                o_ya = 8'd0;
                o_xb = -8'd8;
                o_yb = -8'd4;
            end
            51: begin
                o_xa = 8'd3;
                o_ya = 8'd3;
                o_xb = 8'd7;
                o_yb = 8'd8;
            end
            52: begin
                o_xa = 8'd5;
                o_ya = 8'd7;
                o_xb = 8'd10;
                o_yb = -8'd7;
            end
            53: begin
                o_xa = -8'd1;
                o_ya = 8'd7;
                o_xb = 8'd1;
                o_yb = -8'd12;
            end
            54: begin
                o_xa = 8'd3;
                o_ya = -8'd10;
                o_xb = 8'd5;
                o_yb = 8'd6;
            end
            55: begin
                o_xa = 8'd2;
                o_ya = -8'd4;
                o_xb = 8'd3;
                o_yb = -8'd10;
            end
            56: begin
                o_xa = -8'd13;
                o_ya = 8'd0;
                o_xb = -8'd13;
                o_yb = 8'd5;
            end
            57: begin
                o_xa = -8'd13;
                o_ya = -8'd7;
                o_xb = -8'd12;
                o_yb = 8'd12;
            end
            58: begin
                o_xa = -8'd13;
                o_ya = 8'd3;
                o_xb = -8'd11;
                o_yb = 8'd8;
            end
            59: begin
                o_xa = -8'd7;
                o_ya = 8'd12;
                o_xb = -8'd4;
                o_yb = 8'd7;
            end
            60: begin
                o_xa = 8'd6;
                o_ya = -8'd10;
                o_xb = 8'd12;
                o_yb = 8'd8;
            end
            61: begin
                o_xa = -8'd9;
                o_ya = -8'd1;
                o_xb = -8'd7;
                o_yb = -8'd6;
            end
            62: begin
                o_xa = -8'd2;
                o_ya = -8'd5;
                o_xb = 8'd0;
                o_yb = 8'd12;
            end
            63: begin
                o_xa = -8'd12;
                o_ya = 8'd5;
                o_xb = -8'd7;
                o_yb = 8'd5;
            end
            64: begin
                o_xa = 8'd3;
                o_ya = -8'd10;
                o_xb = 8'd8;
                o_yb = -8'd13;
            end
            65: begin
                o_xa = -8'd7;
                o_ya = -8'd7;
                o_xb = -8'd4;
                o_yb = 8'd5;
            end
            66: begin
                o_xa = -8'd3;
                o_ya = -8'd2;
                o_xb = -8'd1;
                o_yb = -8'd7;
            end
            67: begin
                o_xa = 8'd2;
                o_ya = 8'd9;
                o_xb = 8'd5;
                o_yb = -8'd11;
            end
            68: begin
                o_xa = -8'd11;
                o_ya = -8'd13;
                o_xb = -8'd5;
                o_yb = -8'd13;
            end
            69: begin
                o_xa = -8'd1;
                o_ya = 8'd6;
                o_xb = 8'd0;
                o_yb = -8'd1;
            end
            70: begin
                o_xa = 8'd5;
                o_ya = -8'd3;
                o_xb = 8'd5;
                o_yb = 8'd2;
            end
            71: begin
                o_xa = -8'd4;
                o_ya = -8'd13;
                o_xb = -8'd4;
                o_yb = 8'd12;
            end
            72: begin
                o_xa = -8'd9;
                o_ya = -8'd6;
                o_xb = -8'd9;
                o_yb = 8'd6;
            end
            73: begin
                o_xa = -8'd12;
                o_ya = -8'd10;
                o_xb = -8'd8;
                o_yb = -8'd4;
            end
            74: begin
                o_xa = 8'd10;
                o_ya = 8'd2;
                o_xb = 8'd12;
                o_yb = -8'd3;
            end
            75: begin
                o_xa = 8'd7;
                o_ya = 8'd12;
                o_xb = 8'd12;
                o_yb = 8'd12;
            end
            76: begin
                o_xa = -8'd7;
                o_ya = -8'd13;
                o_xb = -8'd6;
                o_yb = 8'd5;
            end
            77: begin
                o_xa = -8'd4;
                o_ya = 8'd9;
                o_xb = -8'd3;
                o_yb = 8'd4;
            end
            78: begin
                o_xa = 8'd7;
                o_ya = -8'd1;
                o_xb = 8'd12;
                o_yb = 8'd2;
            end
            79: begin
                o_xa = -8'd7;
                o_ya = 8'd6;
                o_xb = -8'd5;
                o_yb = 8'd1;
            end
            80: begin
                o_xa = -8'd13;
                o_ya = 8'd11;
                o_xb = -8'd12;
                o_yb = 8'd5;
            end
            81: begin
                o_xa = -8'd3;
                o_ya = 8'd7;
                o_xb = -8'd2;
                o_yb = -8'd6;
            end
            82: begin
                o_xa = 8'd7;
                o_ya = -8'd8;
                o_xb = 8'd12;
                o_yb = -8'd7;
            end
            83: begin
                o_xa = -8'd13;
                o_ya = -8'd7;
                o_xb = -8'd11;
                o_yb = -8'd12;
            end
            84: begin
                o_xa = 8'd1;
                o_ya = -8'd3;
                o_xb = 8'd12;
                o_yb = 8'd12;
            end
            85: begin
                o_xa = 8'd2;
                o_ya = -8'd6;
                o_xb = 8'd3;
                o_yb = 8'd0;
            end
            86: begin
                o_xa = -8'd4;
                o_ya = 8'd3;
                o_xb = -8'd2;
                o_yb = -8'd13;
            end
            87: begin
                o_xa = -8'd1;
                o_ya = -8'd13;
                o_xb = 8'd1;
                o_yb = 8'd9;
            end
            88: begin
                o_xa = 8'd7;
                o_ya = 8'd1;
                o_xb = 8'd8;
                o_yb = -8'd6;
            end
            89: begin
                o_xa = 8'd1;
                o_ya = -8'd1;
                o_xb = 8'd3;
                o_yb = 8'd12;
            end
            90: begin
                o_xa = 8'd9;
                o_ya = 8'd1;
                o_xb = 8'd12;
                o_yb = 8'd6;
            end
            91: begin
                o_xa = -8'd1;
                o_ya = -8'd9;
                o_xb = -8'd1;
                o_yb = 8'd3;
            end
            92: begin
                o_xa = -8'd13;
                o_ya = -8'd13;
                o_xb = -8'd10;
                o_yb = 8'd5;
            end
            93: begin
                o_xa = 8'd7;
                o_ya = 8'd7;
                o_xb = 8'd10;
                o_yb = 8'd12;
            end
            94: begin
                o_xa = 8'd12;
                o_ya = -8'd5;
                o_xb = 8'd12;
                o_yb = 8'd9;
            end
            95: begin
                o_xa = 8'd6;
                o_ya = 8'd3;
                o_xb = 8'd7;
                o_yb = 8'd11;
            end
            96: begin
                o_xa = 8'd5;
                o_ya = -8'd13;
                o_xb = 8'd6;
                o_yb = 8'd10;
            end
            97: begin
                o_xa = 8'd2;
                o_ya = -8'd12;
                o_xb = 8'd2;
                o_yb = 8'd3;
            end
            98: begin
                o_xa = 8'd3;
                o_ya = 8'd8;
                o_xb = 8'd4;
                o_yb = -8'd6;
            end
            99: begin
                o_xa = 8'd2;
                o_ya = 8'd6;
                o_xb = 8'd12;
                o_yb = -8'd13;
            end
            100: begin
                o_xa = 8'd9;
                o_ya = -8'd12;
                o_xb = 8'd10;
                o_yb = 8'd3;
            end
            101: begin
                o_xa = -8'd8;
                o_ya = 8'd4;
                o_xb = -8'd7;
                o_yb = 8'd9;
            end
            102: begin
                o_xa = -8'd11;
                o_ya = 8'd12;
                o_xb = -8'd4;
                o_yb = -8'd6;
            end
            103: begin
                o_xa = 8'd1;
                o_ya = 8'd12;
                o_xb = 8'd2;
                o_yb = -8'd8;
            end
            104: begin
                o_xa = 8'd6;
                o_ya = -8'd9;
                o_xb = 8'd7;
                o_yb = -8'd4;
            end
            105: begin
                o_xa = 8'd2;
                o_ya = 8'd3;
                o_xb = 8'd3;
                o_yb = -8'd2;
            end
            106: begin
                o_xa = 8'd6;
                o_ya = 8'd3;
                o_xb = 8'd11;
                o_yb = 8'd0;
            end
            107: begin
                o_xa = 8'd3;
                o_ya = -8'd3;
                o_xb = 8'd8;
                o_yb = -8'd8;
            end
            108: begin
                o_xa = 8'd7;
                o_ya = 8'd8;
                o_xb = 8'd9;
                o_yb = 8'd3;
            end
            109: begin
                o_xa = -8'd11;
                o_ya = -8'd5;
                o_xb = -8'd6;
                o_yb = -8'd4;
            end
            110: begin
                o_xa = -8'd10;
                o_ya = 8'd11;
                o_xb = -8'd5;
                o_yb = 8'd10;
            end
            111: begin
                o_xa = -8'd5;
                o_ya = -8'd8;
                o_xb = -8'd3;
                o_yb = 8'd12;
            end
            112: begin
                o_xa = -8'd10;
                o_ya = 8'd5;
                o_xb = -8'd9;
                o_yb = 8'd0;
            end
            113: begin
                o_xa = 8'd8;
                o_ya = -8'd1;
                o_xb = 8'd12;
                o_yb = -8'd6;
            end
            114: begin
                o_xa = 8'd4;
                o_ya = -8'd6;
                o_xb = 8'd6;
                o_yb = -8'd11;
            end
            115: begin
                o_xa = -8'd10;
                o_ya = 8'd12;
                o_xb = -8'd8;
                o_yb = 8'd7;
            end
            116: begin
                o_xa = 8'd4;
                o_ya = -8'd2;
                o_xb = 8'd6;
                o_yb = 8'd7;
            end
            117: begin
                o_xa = -8'd2;
                o_ya = 8'd0;
                o_xb = -8'd2;
                o_yb = 8'd12;
            end
            118: begin
                o_xa = -8'd5;
                o_ya = -8'd8;
                o_xb = -8'd5;
                o_yb = 8'd2;
            end
            119: begin
                o_xa = 8'd7;
                o_ya = -8'd6;
                o_xb = 8'd10;
                o_yb = 8'd12;
            end
            120: begin
                o_xa = -8'd9;
                o_ya = -8'd13;
                o_xb = -8'd8;
                o_yb = -8'd8;
            end
            121: begin
                o_xa = -8'd5;
                o_ya = -8'd13;
                o_xb = -8'd5;
                o_yb = -8'd2;
            end
            122: begin
                o_xa = 8'd8;
                o_ya = -8'd8;
                o_xb = 8'd9;
                o_yb = -8'd13;
            end
            123: begin
                o_xa = -8'd9;
                o_ya = -8'd11;
                o_xb = -8'd9;
                o_yb = 8'd0;
            end
            124: begin
                o_xa = 8'd1;
                o_ya = -8'd8;
                o_xb = 8'd1;
                o_yb = -8'd2;
            end
            125: begin
                o_xa = 8'd7;
                o_ya = -8'd4;
                o_xb = 8'd9;
                o_yb = 8'd1;
            end
            126: begin
                o_xa = -8'd2;
                o_ya = 8'd1;
                o_xb = -8'd1;
                o_yb = -8'd4;
            end
            127: begin
                o_xa = 8'd11;
                o_ya = -8'd6;
                o_xb = 8'd12;
                o_yb = -8'd11;
            end
            128: begin
                o_xa = -8'd12;
                o_ya = -8'd9;
                o_xb = -8'd6;
                o_yb = 8'd4;
            end
            129: begin
                o_xa = 8'd3;
                o_ya = 8'd7;
                o_xb = 8'd7;
                o_yb = 8'd12;
            end
            130: begin
                o_xa = 8'd5;
                o_ya = 8'd5;
                o_xb = 8'd10;
                o_yb = 8'd8;
            end
            131: begin
                o_xa = 8'd0;
                o_ya = -8'd4;
                o_xb = 8'd2;
                o_yb = 8'd8;
            end
            132: begin
                o_xa = -8'd9;
                o_ya = 8'd12;
                o_xb = -8'd5;
                o_yb = -8'd13;
            end
            133: begin
                o_xa = 8'd0;
                o_ya = 8'd7;
                o_xb = 8'd2;
                o_yb = 8'd12;
            end
            134: begin
                o_xa = -8'd1;
                o_ya = 8'd2;
                o_xb = 8'd1;
                o_yb = 8'd7;
            end
            135: begin
                o_xa = 8'd5;
                o_ya = 8'd11;
                o_xb = 8'd7;
                o_yb = -8'd9;
            end
            136: begin
                o_xa = 8'd3;
                o_ya = 8'd5;
                o_xb = 8'd6;
                o_yb = -8'd8;
            end
            137: begin
                o_xa = -8'd13;
                o_ya = -8'd4;
                o_xb = -8'd8;
                o_yb = 8'd9;
            end
            138: begin
                o_xa = -8'd5;
                o_ya = 8'd9;
                o_xb = -8'd3;
                o_yb = -8'd3;
            end
            139: begin
                o_xa = -8'd4;
                o_ya = -8'd7;
                o_xb = -8'd3;
                o_yb = -8'd12;
            end
            140: begin
                o_xa = 8'd6;
                o_ya = 8'd5;
                o_xb = 8'd8;
                o_yb = 8'd0;
            end
            141: begin
                o_xa = -8'd7;
                o_ya = 8'd6;
                o_xb = -8'd6;
                o_yb = 8'd12;
            end
            142: begin
                o_xa = -8'd13;
                o_ya = 8'd6;
                o_xb = -8'd5;
                o_yb = -8'd2;
            end
            143: begin
                o_xa = 8'd1;
                o_ya = -8'd10;
                o_xb = 8'd3;
                o_yb = 8'd10;
            end
            144: begin
                o_xa = 8'd4;
                o_ya = 8'd1;
                o_xb = 8'd8;
                o_yb = -8'd4;
            end
            145: begin
                o_xa = -8'd2;
                o_ya = -8'd2;
                o_xb = 8'd2;
                o_yb = -8'd13;
            end
            146: begin
                o_xa = 8'd2;
                o_ya = -8'd12;
                o_xb = 8'd12;
                o_yb = 8'd12;
            end
            147: begin
                o_xa = -8'd2;
                o_ya = -8'd13;
                o_xb = 8'd0;
                o_yb = -8'd6;
            end
            148: begin
                o_xa = 8'd4;
                o_ya = 8'd1;
                o_xb = 8'd9;
                o_yb = 8'd3;
            end
            149: begin
                o_xa = -8'd6;
                o_ya = -8'd10;
                o_xb = -8'd3;
                o_yb = -8'd5;
            end
            150: begin
                o_xa = -8'd3;
                o_ya = -8'd13;
                o_xb = -8'd1;
                o_yb = 8'd1;
            end
            151: begin
                o_xa = 8'd7;
                o_ya = 8'd5;
                o_xb = 8'd12;
                o_yb = -8'd11;
            end
            152: begin
                o_xa = 8'd4;
                o_ya = -8'd2;
                o_xb = 8'd5;
                o_yb = -8'd7;
            end
            153: begin
                o_xa = -8'd13;
                o_ya = 8'd9;
                o_xb = -8'd9;
                o_yb = -8'd5;
            end
            154: begin
                o_xa = 8'd7;
                o_ya = 8'd1;
                o_xb = 8'd8;
                o_yb = 8'd6;
            end
            155: begin
                o_xa = 8'd7;
                o_ya = -8'd8;
                o_xb = 8'd7;
                o_yb = 8'd6;
            end
            156: begin
                o_xa = -8'd7;
                o_ya = -8'd4;
                o_xb = -8'd7;
                o_yb = 8'd1;
            end
            157: begin
                o_xa = -8'd8;
                o_ya = 8'd11;
                o_xb = -8'd7;
                o_yb = -8'd8;
            end
            158: begin
                o_xa = -8'd13;
                o_ya = 8'd6;
                o_xb = -8'd12;
                o_yb = -8'd8;
            end
            159: begin
                o_xa = 8'd2;
                o_ya = 8'd4;
                o_xb = 8'd3;
                o_yb = 8'd9;
            end
            160: begin
                o_xa = 8'd10;
                o_ya = -8'd5;
                o_xb = 8'd12;
                o_yb = 8'd3;
            end
            161: begin
                o_xa = -8'd6;
                o_ya = -8'd5;
                o_xb = -8'd6;
                o_yb = 8'd7;
            end
            162: begin
                o_xa = 8'd8;
                o_ya = -8'd3;
                o_xb = 8'd9;
                o_yb = -8'd8;
            end
            163: begin
                o_xa = 8'd2;
                o_ya = -8'd12;
                o_xb = 8'd2;
                o_yb = 8'd8;
            end
            164: begin
                o_xa = -8'd11;
                o_ya = -8'd2;
                o_xb = -8'd10;
                o_yb = 8'd3;
            end
            165: begin
                o_xa = -8'd12;
                o_ya = -8'd13;
                o_xb = -8'd7;
                o_yb = -8'd9;
            end
            166: begin
                o_xa = -8'd11;
                o_ya = 8'd0;
                o_xb = -8'd10;
                o_yb = -8'd5;
            end
            167: begin
                o_xa = 8'd5;
                o_ya = -8'd3;
                o_xb = 8'd11;
                o_yb = 8'd8;
            end
            168: begin
                o_xa = -8'd2;
                o_ya = -8'd13;
                o_xb = -8'd1;
                o_yb = 8'd12;
            end
            169: begin
                o_xa = -8'd1;
                o_ya = -8'd8;
                o_xb = 8'd0;
                o_yb = 8'd9;
            end
            170: begin
                o_xa = -8'd13;
                o_ya = -8'd11;
                o_xb = -8'd12;
                o_yb = -8'd5;
            end
            171: begin
                o_xa = -8'd10;
                o_ya = -8'd2;
                o_xb = -8'd10;
                o_yb = 8'd11;
            end
            172: begin
                o_xa = -8'd3;
                o_ya = 8'd9;
                o_xb = -8'd2;
                o_yb = -8'd13;
            end
            173: begin
                o_xa = 8'd2;
                o_ya = -8'd3;
                o_xb = 8'd3;
                o_yb = 8'd2;
            end
            174: begin
                o_xa = -8'd9;
                o_ya = -8'd13;
                o_xb = -8'd4;
                o_yb = 8'd0;
            end
            175: begin
                o_xa = -8'd4;
                o_ya = 8'd6;
                o_xb = -8'd3;
                o_yb = -8'd10;
            end
            176: begin
                o_xa = -8'd4;
                o_ya = 8'd12;
                o_xb = -8'd2;
                o_yb = -8'd7;
            end
            177: begin
                o_xa = -8'd6;
                o_ya = -8'd11;
                o_xb = -8'd4;
                o_yb = 8'd9;
            end
            178: begin
                o_xa = 8'd6;
                o_ya = -8'd3;
                o_xb = 8'd6;
                o_yb = 8'd11;
            end
            179: begin
                o_xa = -8'd13;
                o_ya = 8'd11;
                o_xb = -8'd5;
                o_yb = 8'd5;
            end
            180: begin
                o_xa = 8'd11;
                o_ya = 8'd11;
                o_xb = 8'd12;
                o_yb = 8'd6;
            end
            181: begin
                o_xa = 8'd7;
                o_ya = -8'd5;
                o_xb = 8'd12;
                o_yb = -8'd2;
            end
            182: begin
                o_xa = -8'd1;
                o_ya = 8'd12;
                o_xb = 8'd0;
                o_yb = 8'd7;
            end
            183: begin
                o_xa = -8'd4;
                o_ya = -8'd8;
                o_xb = -8'd3;
                o_yb = -8'd2;
            end
            184: begin
                o_xa = -8'd7;
                o_ya = 8'd1;
                o_xb = -8'd6;
                o_yb = 8'd7;
            end
            185: begin
                o_xa = -8'd13;
                o_ya = -8'd12;
                o_xb = -8'd8;
                o_yb = -8'd13;
            end
            186: begin
                o_xa = -8'd7;
                o_ya = -8'd2;
                o_xb = -8'd6;
                o_yb = -8'd8;
            end
            187: begin
                o_xa = -8'd8;
                o_ya = 8'd5;
                o_xb = -8'd6;
                o_yb = -8'd9;
            end
            188: begin
                o_xa = -8'd5;
                o_ya = -8'd1;
                o_xb = -8'd4;
                o_yb = 8'd5;
            end
            189: begin
                o_xa = -8'd13;
                o_ya = 8'd7;
                o_xb = -8'd8;
                o_yb = 8'd10;
            end
            190: begin
                o_xa = 8'd1;
                o_ya = 8'd5;
                o_xb = 8'd5;
                o_yb = -8'd13;
            end
            191: begin
                o_xa = 8'd1;
                o_ya = 8'd0;
                o_xb = 8'd10;
                o_yb = -8'd13;
            end
            192: begin
                o_xa = 8'd9;
                o_ya = 8'd12;
                o_xb = 8'd10;
                o_yb = -8'd1;
            end
            193: begin
                o_xa = 8'd5;
                o_ya = -8'd8;
                o_xb = 8'd10;
                o_yb = -8'd9;
            end
            194: begin
                o_xa = -8'd1;
                o_ya = 8'd11;
                o_xb = 8'd1;
                o_yb = -8'd13;
            end
            195: begin
                o_xa = -8'd9;
                o_ya = -8'd3;
                o_xb = -8'd6;
                o_yb = 8'd2;
            end
            196: begin
                o_xa = -8'd1;
                o_ya = -8'd10;
                o_xb = 8'd1;
                o_yb = 8'd12;
            end
            197: begin
                o_xa = -8'd13;
                o_ya = 8'd1;
                o_xb = -8'd8;
                o_yb = -8'd10;
            end
            198: begin
                o_xa = 8'd8;
                o_ya = -8'd11;
                o_xb = 8'd10;
                o_yb = -8'd6;
            end
            199: begin
                o_xa = 8'd2;
                o_ya = -8'd13;
                o_xb = 8'd3;
                o_yb = -8'd6;
            end
            200: begin
                o_xa = 8'd7;
                o_ya = -8'd13;
                o_xb = 8'd12;
                o_yb = -8'd9;
            end
            201: begin
                o_xa = -8'd10;
                o_ya = -8'd10;
                o_xb = -8'd5;
                o_yb = -8'd7;
            end
            202: begin
                o_xa = -8'd10;
                o_ya = -8'd8;
                o_xb = -8'd8;
                o_yb = -8'd13;
            end
            203: begin
                o_xa = 8'd4;
                o_ya = -8'd6;
                o_xb = 8'd8;
                o_yb = 8'd5;
            end
            204: begin
                o_xa = 8'd3;
                o_ya = 8'd12;
                o_xb = 8'd8;
                o_yb = -8'd13;
            end
            205: begin
                o_xa = -8'd4;
                o_ya = 8'd2;
                o_xb = -8'd3;
                o_yb = -8'd3;
            end
            206: begin
                o_xa = 8'd5;
                o_ya = -8'd13;
                o_xb = 8'd10;
                o_yb = -8'd12;
            end
            207: begin
                o_xa = 8'd4;
                o_ya = -8'd13;
                o_xb = 8'd5;
                o_yb = -8'd1;
            end
            208: begin
                o_xa = -8'd9;
                o_ya = 8'd9;
                o_xb = -8'd4;
                o_yb = 8'd3;
            end
            209: begin
                o_xa = 8'd0;
                o_ya = 8'd3;
                o_xb = 8'd3;
                o_yb = -8'd9;
            end
            210: begin
                o_xa = -8'd12;
                o_ya = 8'd1;
                o_xb = -8'd6;
                o_yb = 8'd1;
            end
            211: begin
                o_xa = 8'd3;
                o_ya = 8'd2;
                o_xb = 8'd4;
                o_yb = -8'd8;
            end
            212: begin
                o_xa = -8'd10;
                o_ya = -8'd10;
                o_xb = -8'd10;
                o_yb = 8'd9;
            end
            213: begin
                o_xa = 8'd8;
                o_ya = -8'd13;
                o_xb = 8'd12;
                o_yb = 8'd12;
            end
            214: begin
                o_xa = -8'd8;
                o_ya = -8'd12;
                o_xb = -8'd6;
                o_yb = -8'd5;
            end
            215: begin
                o_xa = 8'd2;
                o_ya = 8'd2;
                o_xb = 8'd3;
                o_yb = 8'd7;
            end
            216: begin
                o_xa = 8'd10;
                o_ya = 8'd6;
                o_xb = 8'd11;
                o_yb = -8'd8;
            end
            217: begin
                o_xa = 8'd6;
                o_ya = 8'd8;
                o_xb = 8'd8;
                o_yb = -8'd12;
            end
            218: begin
                o_xa = -8'd7;
                o_ya = 8'd10;
                o_xb = -8'd6;
                o_yb = 8'd5;
            end
            219: begin
                o_xa = -8'd3;
                o_ya = -8'd9;
                o_xb = -8'd3;
                o_yb = 8'd9;
            end
            220: begin
                o_xa = -8'd1;
                o_ya = -8'd13;
                o_xb = -8'd1;
                o_yb = 8'd5;
            end
            221: begin
                o_xa = -8'd3;
                o_ya = -8'd7;
                o_xb = -8'd3;
                o_yb = 8'd4;
            end
            222: begin
                o_xa = -8'd8;
                o_ya = -8'd2;
                o_xb = -8'd8;
                o_yb = 8'd3;
            end
            223: begin
                o_xa = 8'd4;
                o_ya = 8'd2;
                o_xb = 8'd12;
                o_yb = 8'd12;
            end
            224: begin
                o_xa = 8'd2;
                o_ya = -8'd5;
                o_xb = 8'd3;
                o_yb = 8'd11;
            end
            225: begin
                o_xa = 8'd6;
                o_ya = -8'd9;
                o_xb = 8'd11;
                o_yb = -8'd13;
            end
            226: begin
                o_xa = 8'd3;
                o_ya = -8'd1;
                o_xb = 8'd7;
                o_yb = 8'd12;
            end
            227: begin
                o_xa = 8'd11;
                o_ya = -8'd1;
                o_xb = 8'd12;
                o_yb = 8'd4;
            end
            228: begin
                o_xa = -8'd3;
                o_ya = 8'd0;
                o_xb = -8'd3;
                o_yb = 8'd6;
            end
            229: begin
                o_xa = 8'd4;
                o_ya = -8'd11;
                o_xb = 8'd4;
                o_yb = 8'd12;
            end
            230: begin
                o_xa = 8'd2;
                o_ya = -8'd4;
                o_xb = 8'd2;
                o_yb = 8'd1;
            end
            231: begin
                o_xa = -8'd10;
                o_ya = -8'd6;
                o_xb = -8'd8;
                o_yb = 8'd1;
            end
            232: begin
                o_xa = -8'd13;
                o_ya = 8'd7;
                o_xb = -8'd11;
                o_yb = 8'd1;
            end
            233: begin
                o_xa = -8'd13;
                o_ya = 8'd12;
                o_xb = -8'd11;
                o_yb = -8'd13;
            end
            234: begin
                o_xa = 8'd6;
                o_ya = 8'd0;
                o_xb = 8'd11;
                o_yb = -8'd13;
            end
            235: begin
                o_xa = 8'd0;
                o_ya = -8'd1;
                o_xb = 8'd1;
                o_yb = 8'd4;
            end
            236: begin
                o_xa = -8'd13;
                o_ya = 8'd3;
                o_xb = -8'd9;
                o_yb = -8'd2;
            end
            237: begin
                o_xa = -8'd9;
                o_ya = 8'd8;
                o_xb = -8'd6;
                o_yb = -8'd3;
            end
            238: begin
                o_xa = -8'd13;
                o_ya = -8'd6;
                o_xb = -8'd8;
                o_yb = -8'd2;
            end
            239: begin
                o_xa = 8'd5;
                o_ya = -8'd9;
                o_xb = 8'd8;
                o_yb = 8'd10;
            end
            240: begin
                o_xa = 8'd2;
                o_ya = 8'd7;
                o_xb = 8'd3;
                o_yb = -8'd9;
            end
            241: begin
                o_xa = -8'd1;
                o_ya = -8'd6;
                o_xb = -8'd1;
                o_yb = -8'd1;
            end
            242: begin
                o_xa = 8'd9;
                o_ya = 8'd5;
                o_xb = 8'd11;
                o_yb = -8'd2;
            end
            243: begin
                o_xa = 8'd11;
                o_ya = -8'd3;
                o_xb = 8'd12;
                o_yb = -8'd8;
            end
            244: begin
                o_xa = 8'd3;
                o_ya = 8'd0;
                o_xb = 8'd3;
                o_yb = 8'd5;
            end
            245: begin
                o_xa = -8'd1;
                o_ya = 8'd4;
                o_xb = 8'd0;
                o_yb = 8'd10;
            end
            246: begin
                o_xa = 8'd3;
                o_ya = -8'd6;
                o_xb = 8'd4;
                o_yb = 8'd5;
            end
            247: begin
                o_xa = -8'd13;
                o_ya = 8'd0;
                o_xb = -8'd10;
                o_yb = 8'd5;
            end
            248: begin
                o_xa = 8'd5;
                o_ya = 8'd8;
                o_xb = 8'd12;
                o_yb = 8'd11;
            end
            249: begin
                o_xa = 8'd8;
                o_ya = 8'd9;
                o_xb = 8'd9;
                o_yb = -8'd6;
            end
            250: begin
                o_xa = 8'd7;
                o_ya = -8'd4;
                o_xb = 8'd8;
                o_yb = -8'd12;
            end
            251: begin
                o_xa = -8'd10;
                o_ya = 8'd4;
                o_xb = -8'd10;
                o_yb = 8'd9;
            end
            252: begin
                o_xa = 8'd7;
                o_ya = 8'd3;
                o_xb = 8'd12;
                o_yb = 8'd4;
            end
            253: begin
                o_xa = 8'd9;
                o_ya = -8'd7;
                o_xb = 8'd10;
                o_yb = -8'd2;
            end
            254: begin
                o_xa = 8'd7;
                o_ya = 8'd0;
                o_xb = 8'd12;
                o_yb = -8'd2;
            end
            255: begin
                o_xa = -8'd1;
                o_ya = -8'd6;
                o_xb = 8'd0;
                o_yb = -8'd11;
            end
        endcase
    end
endmodule