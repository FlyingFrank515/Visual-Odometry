`include "MATCH.v"
`include "Key_Buffer2.v"

module MATCH_Top
#(
    
)
(

)
endmodule
